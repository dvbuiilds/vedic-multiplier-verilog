//: version "2.1"
//: property encoding = "utf-8"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "BIN-TO-BCD.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg w0;    //: /sn:0 {0}(73,66)(73,92){1}
//: {2}(75,94)(91,94)(91,109){3}
//: {4}(73,96)(73,154){5}
//: {6}(75,156)(85,156)(85,155)(433,155){7}
//: {8}(73,158)(73,186){9}
//: {10}(75,188)(85,188)(85,190)(433,190){11}
//: {12}(73,190)(73,235){13}
//: {14}(75,237)(85,237)(85,236)(457,236){15}
//: {16}(73,239)(73,346){17}
//: {18}(75,348)(85,348)(85,349)(400,349){19}
//: {20}(73,350)(73,473){21}
reg w3;    //: /sn:0 {0}(359,64)(359,441)(560,441){1}
reg w1;    //: /sn:0 {0}(432,285)(179,285){1}
//: {2}(177,283)(177,162){3}
//: {4}(179,160)(433,160){5}
//: {6}(177,158)(177,93){7}
//: {8}(179,91)(194,91)(194,110){9}
//: {10}(177,89)(177,65){11}
//: {12}(177,287)(177,315){13}
//: {14}(179,317)(189,317)(189,315)(433,315){15}
//: {16}(177,319)(177,354){17}
//: {18}(179,356)(189,356)(189,354)(400,354){19}
//: {20}(177,358)(177,468){21}
reg w2;    //: /sn:0 {0}(433,320)(271,320){1}
//: {2}(269,318)(269,196){3}
//: {4}(271,194)(281,194)(281,195)(433,195){5}
//: {6}(269,192)(269,97){7}
//: {8}(271,95)(281,95)(281,101)(288,101)(288,111){9}
//: {10}(269,93)(269,64){11}
//: {12}(269,322)(269,394){13}
//: {14}(271,396)(432,396){15}
//: {16}(269,398)(269,470){17}
wire w7;    //: /sn:0 {0}(194,126)(194,241){1}
//: {2}(196,243)(206,243)(206,246)(399,246){3}
//: {4}(194,245)(194,470){5}
wire w34;    //: /sn:0 {0}(454,193)(481,193)(481,177)(496,177){1}
wire w39;    //: /sn:0 {0}(472,363)(485,363)(485,377)(500,377){1}
wire w36;    //: /sn:0 {0}(453,283)(483,283)(483,299)(498,299){1}
wire w20;    //: /sn:0 {0}(478,239)(556,239){1}
wire w30;    //: /sn:0 {0}(91,125)(91,277){1}
//: {2}(93,279)(103,279)(103,280)(432,280){3}
//: {4}(91,281)(91,385){5}
//: {6}(93,387)(103,387)(103,391)(432,391){7}
//: {8}(91,389)(91,473){9}
wire w37;    //: /sn:0 {0}(454,318)(483,318)(483,304)(498,304){1}
wire w19;    //: /sn:0 {0}(420,249)(442,249)(442,241)(457,241){1}
wire w32;    //: /sn:0 {0}(453,394)(485,394)(485,382)(500,382){1}
wire w27;    //: /sn:0 {0}(421,352)(436,352)(436,360)(451,360){1}
wire w28;    //: /sn:0 {0}(288,127)(288,249){1}
//: {2}(290,251)(399,251){3}
//: {4}(288,253)(288,364){5}
//: {6}(290,366)(300,366)(300,365)(451,365){7}
//: {8}(288,368)(288,469){9}
wire w33;    //: /sn:0 {0}(454,158)(481,158)(481,172)(496,172){1}
wire w35;    //: /sn:0 {0}(517,175)(557,175){1}
wire w41;    //: /sn:0 {0}(521,380)(562,380){1}
wire w38;    //: /sn:0 {0}(519,302)(559,302){1}
//: enddecls

  //: comment g44 @(175,7) /sn:0
  //: /line:"B"
  //: /end
  _GGNBUF #(2) g4 (.I(w0), .Z(w30));   //: @(91,115) /sn:0 /R:3 /w:[ 3 0 ]
  _GGAND2 #(6) g8 (.I0(w0), .I1(w1), .Z(w33));   //: @(444,158) /sn:0 /w:[ 7 5 0 ]
  //: comment g47 @(605,165) /sn:0
  //: /line:"B5"
  //: /end
  //: SWITCH g3 (w3) @(359,51) /sn:0 /R:3 /w:[ 0 ] /st:0 /dn:1
  _GGOR2 #(6) g16 (.I0(w36), .I1(w37), .Z(w38));   //: @(509,302) /sn:0 /w:[ 1 1 0 ]
  //: joint g26 (w0) @(73, 348) /w:[ 18 17 -1 20 ]
  _GGOR2 #(6) g17 (.I0(w39), .I1(w32), .Z(w41));   //: @(511,380) /sn:0 /w:[ 1 1 0 ]
  //: SWITCH g2 (w2) @(269,51) /sn:0 /R:3 /w:[ 11 ] /st:0 /dn:1
  //: joint g30 (w30) @(91, 279) /w:[ 2 1 -1 4 ]
  //: joint g23 (w2) @(269, 396) /w:[ 14 13 -1 16 ]
  //: LED g39 (w20) @(563,239) /sn:0 /R:3 /w:[ 1 ] /type:0
  //: joint g24 (w30) @(91, 387) /w:[ 6 5 -1 8 ]
  //: SWITCH g1 (w1) @(177,52) /sn:0 /R:3 /w:[ 11 ] /st:0 /dn:1
  //: joint g29 (w1) @(177, 285) /w:[ 1 2 -1 12 ]
  //: comment g51 @(604,434) /sn:0
  //: /line:"B5"
  //: /end
  _GGAND2 #(6) g18 (.I0(w0), .I1(w1), .Z(w27));   //: @(411,352) /sn:0 /w:[ 19 19 0 ]
  //: joint g25 (w1) @(177, 356) /w:[ 18 17 -1 20 ]
  _GGAND2 #(6) g10 (.I0(w0), .I1(w19), .Z(w20));   //: @(468,239) /sn:0 /w:[ 15 1 0 ]
  //: comment g49 @(605,298) /sn:0
  //: /line:"B3"
  //: /end
  //: comment g50 @(603,374) /sn:0
  //: /line:"B4"
  //: /end
  _GGNBUF #(2) g6 (.I(w2), .Z(w28));   //: @(288,117) /sn:0 /R:3 /w:[ 9 0 ]
  //: joint g35 (w0) @(73, 188) /w:[ 10 9 -1 12 ]
  _GGAND2 #(6) g7 (.I0(w7), .I1(w28), .Z(w19));   //: @(410,249) /sn:0 /w:[ 3 3 0 ]
  _GGAND2 #(6) g9 (.I0(w0), .I1(w2), .Z(w34));   //: @(444,193) /sn:0 /w:[ 11 5 0 ]
  //: joint g31 (w28) @(288, 251) /w:[ 2 1 -1 4 ]
  //: joint g22 (w28) @(288, 366) /w:[ 6 5 -1 8 ]
  //: comment g45 @(265,5) /sn:0
  //: /line:"C"
  //: /end
  //: LED g41 (w41) @(569,380) /sn:0 /R:3 /w:[ 1 ] /type:0
  //: joint g36 (w1) @(177, 160) /w:[ 4 6 -1 3 ]
  //: joint g33 (w0) @(73, 237) /w:[ 14 13 -1 16 ]
  //: LED g42 (w3) @(567,441) /sn:0 /R:3 /w:[ 1 ] /type:0
  //: LED g40 (w38) @(566,302) /sn:0 /R:3 /w:[ 1 ] /type:0
  _GGAND2 #(6) g12 (.I0(w1), .I1(w2), .Z(w37));   //: @(444,318) /sn:0 /w:[ 15 0 0 ]
  //: comment g46 @(355,9) /sn:0
  //: /line:"D"
  //: /end
  //: joint g34 (w2) @(269, 194) /w:[ 4 6 -1 3 ]
  //: joint g28 (w2) @(269, 320) /w:[ 1 2 -1 12 ]
  _GGNBUF #(2) g5 (.I(w1), .Z(w7));   //: @(194,116) /sn:0 /R:3 /w:[ 9 0 ]
  _GGAND2 #(6) g11 (.I0(w30), .I1(w1), .Z(w36));   //: @(443,283) /sn:0 /w:[ 3 0 0 ]
  _GGAND2 #(6) g14 (.I0(w30), .I1(w2), .Z(w32));   //: @(443,394) /sn:0 /w:[ 7 15 0 ]
  //: joint g21 (w0) @(73, 94) /w:[ 2 1 -1 4 ]
  //: joint g19 (w2) @(269, 95) /w:[ 8 10 -1 7 ]
  //: joint g32 (w7) @(194, 243) /w:[ 2 1 -1 4 ]
  //: joint g20 (w1) @(177, 91) /w:[ 8 10 -1 7 ]
  //: comment g43 @(62,7) /sn:0
  //: /line:"A"
  //: /line:""
  //: /end
  //: LED g38 (w35) @(564,175) /sn:0 /R:3 /w:[ 1 ] /type:0
  //: SWITCH g0 (w0) @(73,53) /sn:0 /R:3 /w:[ 0 ] /st:1 /dn:1
  _GGOR2 #(6) g15 (.I0(w33), .I1(w34), .Z(w35));   //: @(507,175) /sn:0 /w:[ 1 1 0 ]
  //: comment g48 @(605,230) /sn:0
  //: /line:"B4"
  //: /end
  //: joint g27 (w1) @(177, 317) /w:[ 14 13 -1 16 ]
  //: joint g37 (w0) @(73, 156) /w:[ 6 5 -1 8 ]
  _GGAND2 #(6) g13 (.I0(w27), .I1(w28), .Z(w39));   //: @(462,363) /sn:0 /w:[ 1 7 0 ]

endmodule
//: /netlistEnd

