//: version "2.1"
//: property encoding = "utf-8"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "new.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg w6;    //: /sn:0 {0}(214,270)(214,115)(291,115){1}
//: {2}(295,115)(383,115){3}
//: {4}(387,115)(447,115){5}
//: {6}(451,115)(454,115)(454,214)(810,214)(810,299){7}
//: {8}(449,113)(449,103)(594,103)(594,400){9}
//: {10}(385,117)(385,319){11}
//: {12}(293,113)(293,100){13}
reg w7;    //: /sn:0 {0}(95,290)(95,153)(112,153){1}
//: {2}(114,151)(114,131){3}
//: {4}(116,129)(238,129){5}
//: {6}(242,129)(626,129)(626,400){7}
//: {8}(240,131)(240,214)(337,214)(337,319){9}
//: {10}(114,127)(114,99){11}
//: {12}(114,155)(114,223)(182,223)(182,270){13}
reg w4;    //: /sn:0 {0}(915,279)(915,201)(779,201){1}
//: {2}(775,201)(665,201){3}
//: {4}(663,199)(663,102){5}
//: {6}(661,201)(580,201){7}
//: {8}(576,201)(417,201)(417,319){9}
//: {10}(578,203)(578,400){11}
//: {12}(777,203)(777,213)(778,213)(778,299){13}
reg w3;    //: /sn:0 {0}(931,279)(931,192)(795,192){1}
//: {2}(791,192)(718,192){3}
//: {4}(716,190)(716,173){5}
//: {6}(714,192)(612,192){7}
//: {8}(608,192)(572,192)(572,180)(353,180)(353,319){9}
//: {10}(610,194)(610,400){11}
//: {12}(793,194)(793,204)(794,204)(794,299){13}
reg w0;    //: /sn:0 {0}(100,290)(100,196)(153,196){1}
//: {2}(157,196)(166,196)(166,270){3}
//: {4}(155,194)(155,184)(170,184)(170,195)(155,195)(155,186){5}
//: {6}(155,198)(155,203)(399,203){7}
//: {8}(403,203)(411,203)(411,256)(530,256)(530,400){9}
//: {10}(401,205)(401,319){11}
reg w1;    //: /sn:0 {0}(198,270)(198,193)(334,193){1}
//: {2}(338,193)(365,193){3}
//: {4}(369,193)(515,193){5}
//: {6}(519,193)(562,193)(562,400){7}
//: {8}(517,195)(517,224)(746,224)(746,299){9}
//: {10}(367,195)(367,253)(369,253)(369,319){11}
//: {12}(336,191)(336,178){13}
reg w2;    //: /sn:0 {0}(642,400)(642,182)(824,182){1}
//: {2}(828,182)(916,182){3}
//: {4}(920,182)(961,182){5}
//: {6}(965,182)(1008,182)(1008,282){7}
//: {8}(963,184)(963,279){9}
//: {10}(918,180)(918,176){11}
//: {12}(826,184)(826,299){13}
reg w5;    //: /sn:0 {0}(855,100)(855,121){1}
//: {2}(857,123)(945,123){3}
//: {4}(949,123)(1013,123)(1013,282){5}
//: {6}(947,125)(947,279){7}
//: {8}(853,123)(762,123)(762,124){9}
//: {10}(760,126)(546,126)(546,400){11}
//: {12}(762,128)(762,299){13}
wire w16;    //: /sn:0 {0}(129,638)(129,702)(186,702)(186,720){1}
wire w13;    //: /sn:0 {0}(97,311)(97,525){1}
wire w34;    //: /sn:0 {0}(756,671)(756,685)(690,685)(690,544)(570,544)(570,559){1}
wire w25;    //: /sn:0 {0}(642,501)(642,528)(740,528)(740,558){1}
wire w22;    //: /sn:0 {0}(401,426)(401,524)(243,524)(243,571){1}
wire w20;    //: /sn:0 {0}(810,406)(810,528)(756,528)(756,558){1}
wire w30;    //: /sn:0 {0}(899,642)(899,650)(850,650)(850,541)(772,541)(772,558){1}
wire w29;    //: /sn:0 {0}(259,684)(259,700)(313,700)(313,715){1}
wire w42;    //: /sn:0 {0}(915,642)(915,702)(891,702)(891,717){1}
wire w12;    //: /sn:0 {0}(113,718)(113,638){1}
wire w19;    //: /sn:0 {0}(963,374)(963,711){1}
wire w18;    //: /sn:0 {0}(947,374)(947,511)(915,511)(915,541){1}
wire w23;    //: /sn:0 {0}(417,426)(417,529)(538,529)(538,559){1}
wire w10;    //: /sn:0 {0}(1010,303)(1010,713){1}
wire w24;    //: /sn:0 {0}(626,501)(626,529)(554,529)(554,559){1}
wire w21;    //: /sn:0 {0}(826,406)(826,443)(899,443)(899,541){1}
wire w27;    //: /sn:0 {0}(554,672)(554,681)(467,681)(467,556)(259,556)(259,571){1}
wire w33;    //: /sn:0 {0}(772,671)(772,705)(748,705)(748,720){1}
wire w14;    //: /sn:0 {0}(198,365)(198,485)(113,485)(113,525){1}
wire w11;    //: /sn:0 {0}(243,684)(243,691)(190,691)(190,517)(129,517)(129,525){1}
wire w15;    //: /sn:0 {0}(214,365)(214,541)(227,541)(227,571){1}
wire w38;    //: /sn:0 {0}(554,716)(554,697)(570,697)(570,672){1}
//: enddecls

  //: LED g44 (w12) @(113,725) /sn:0 /R:2 /w:[ 0 ] /type:0
  _GGAND2 #(6) g8 (.I0(w5), .I1(w2), .Z(w10));   //: @(1010,293) /sn:0 /R:3 /w:[ 5 7 0 ]
  //: SWITCH g4 (w4) @(663,89) /sn:0 /R:3 /w:[ 5 ] /st:1 /dn:0
  //: LED g47 (w38) @(554,723) /sn:0 /R:2 /w:[ 0 ] /type:0
  cross_three g16 (.w0(w2), .w1(w6), .w2(w3), .w3(w4), .w4(w5), .w5(w1), .w6(w21), .w7(w20));   //: @(730, 300) /sz:(112, 105) /R:3 /sn:0 /p:[ Ti0>13 Ti1>7 Ti2>13 Ti3>13 Ti4>13 Ti5>9 Bo0<0 Bo1<0 ]
  //: SWITCH g3 (w3) @(716,160) /sn:0 /R:3 /w:[ 5 ] /st:1 /dn:0
  //: joint g26 (w6) @(449, 115) /w:[ 6 8 5 -1 ]
  //: joint g17 (w2) @(918, 182) /w:[ 4 10 3 -1 ]
  //: SWITCH g2 (w2) @(918,163) /sn:0 /R:3 /w:[ 11 ] /st:0 /dn:0
  //: joint g30 (w5) @(762, 126) /w:[ -1 9 10 12 ]
  cross_four g23 (.w0(w2), .w1(w7), .w2(w3), .w3(w6), .w4(w4), .w5(w1), .w6(w5), .w7(w0), .w8(w25), .w9(w24));   //: @(514, 401) /sz:(144, 99) /R:3 /sn:0 /p:[ Ti0>0 Ti1>7 Ti2>11 Ti3>9 Ti4>11 Ti5>7 Ti6>11 Ti7>9 Bo0<0 Bo1<0 ]
  full_adder g39 (.w8(w27), .w9(w22), .w10(w15), .w0(w29), .w1(w11));   //: @(211, 572) /sz:(64, 111) /R:3 /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Bo0<0 Bo1<0 ]
  //: joint g24 (w2) @(826, 182) /w:[ 2 -1 1 12 ]
  //: SWITCH g1 (w1) @(336,165) /sn:0 /R:3 /w:[ 13 ] /st:1 /dn:0
  //: joint g29 (w1) @(517, 193) /w:[ 6 -1 5 8 ]
  //: LED g51 (w33) @(748,727) /sn:0 /R:2 /w:[ 1 ] /type:0
  //: joint g18 (w6) @(293, 115) /w:[ 2 12 1 -1 ]
  //: joint g25 (w7) @(114, 129) /w:[ 4 10 -1 3 ]
  cross_two g10 (.w0(w2), .w1(w5), .w2(w3), .w3(w4), .w4(w19), .w5(w18));   //: @(899, 280) /sz:(80, 93) /R:3 /sn:0 /p:[ Ti0>9 Ti1>7 Ti2>0 Ti3>0 Bo0<0 Bo1<0 ]
  //: LED g49 (w42) @(891,724) /sn:0 /R:2 /w:[ 1 ] /type:0
  //: LED g50 (w10) @(1010,720) /sn:0 /R:2 /w:[ 1 ] /type:0
  //: SWITCH g6 (w6) @(293,87) /sn:0 /R:3 /w:[ 13 ] /st:0 /dn:0
  //: joint g35 (w6) @(385, 115) /w:[ 4 -1 3 10 ]
  _GGAND2 #(6) g9 (.I0(w0), .I1(w7), .Z(w13));   //: @(97,301) /sn:0 /R:3 /w:[ 0 0 0 ]
  //: SWITCH g7 (w7) @(114,86) /sn:0 /R:3 /w:[ 11 ] /st:1 /dn:0
  cross_three g31 (.w0(w4), .w1(w0), .w2(w6), .w3(w1), .w4(w3), .w5(w7), .w6(w23), .w7(w22));   //: @(321, 320) /sz:(112, 105) /R:3 /sn:0 /p:[ Ti0>9 Ti1>11 Ti2>11 Ti3>11 Ti4>9 Ti5>9 Bo0<0 Bo1<0 ]
  //: joint g22 (w1) @(336, 193) /w:[ 2 12 1 -1 ]
  //: LED g45 (w19) @(963,718) /sn:0 /R:2 /w:[ 1 ] /type:0
  full_adder g41 (.w8(w30), .w9(w20), .w10(w25), .w0(w33), .w1(w34));   //: @(724, 559) /sz:(64, 111) /R:3 /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Bo0<0 Bo1<0 ]
  //: joint g36 (w0) @(401, 203) /w:[ 8 -1 7 10 ]
  //: joint g33 (w3) @(610, 192) /w:[ 7 -1 8 10 ]
  //: comment g52 @(109,54) /sn:0
  //: /line:"a3                             a2                                                         a1                               a0"
  //: /end
  half_adder g40 (.w1(w21), .w0(w18), .w5(w30), .w4(w42));   //: @(883, 542) /sz:(48, 99) /R:3 /sn:0 /p:[ Ti0>1 Ti1>1 Bo0<0 Bo1<0 ]
  full_adder g42 (.w8(w34), .w9(w24), .w10(w23), .w0(w38), .w1(w27));   //: @(522, 560) /sz:(64, 111) /R:3 /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Bo0<1 Bo1<0 ]
  //: joint g12 (w2) @(963, 182) /w:[ 6 -1 5 8 ]
  //: LED g46 (w29) @(313,722) /sn:0 /R:2 /w:[ 1 ] /type:0
  //: joint g34 (w1) @(367, 193) /w:[ 4 -1 3 10 ]
  //: joint g28 (w4) @(663, 201) /w:[ 3 4 6 -1 ]
  //: joint g14 (w0) @(155, 196) /w:[ 2 4 1 6 ]
  //: joint g11 (w5) @(947, 123) /w:[ 4 -1 3 6 ]
  //: SWITCH g5 (w5) @(855,87) /sn:0 /R:3 /w:[ 0 ] /st:0 /dn:0
  //: joint g21 (w5) @(855, 123) /w:[ 2 1 8 -1 ]
  //: joint g19 (w3) @(793, 192) /w:[ 1 -1 2 12 ]
  //: joint g32 (w7) @(240, 129) /w:[ 6 -1 5 8 ]
  //: joint g20 (w4) @(777, 201) /w:[ 1 -1 2 12 ]
  //: LED g43 (w16) @(186,727) /sn:0 /R:2 /w:[ 1 ] /type:0
  full_adder g38 (.w8(w11), .w9(w14), .w10(w13), .w0(w16), .w1(w12));   //: @(81, 526) /sz:(64, 111) /R:3 /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Bo0<0 Bo1<1 ]
  //: joint g15 (w7) @(114, 153) /w:[ -1 2 1 12 ]
  //: SWITCH g0 (w0) @(155,173) /sn:0 /R:3 /w:[ 5 ] /st:0 /dn:0
  //: comment g48 @(111,740) /sn:0
  //: /line:"p7          p6                    p5                                      p4                            p3                       p2          p1      p0"
  //: /end
  //: joint g27 (w3) @(716, 192) /w:[ 3 4 6 -1 ]
  //: joint g37 (w4) @(578, 201) /w:[ 7 -1 8 10 ]
  //: comment g53 @(147,131) /sn:0
  //: /line:"b3                             b2                                                              b1                               b0"
  //: /end
  cross_two g13 (.w0(w6), .w1(w1), .w2(w7), .w3(w0), .w4(w15), .w5(w14));   //: @(150, 271) /sz:(80, 93) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>13 Ti3>3 Bo0<0 Bo1<0 ]

endmodule
//: /netlistEnd

//: /netlistBegin half_adder
module half_adder(w5, w4, w1, w0);
//: interface  /sz:(99, 48) /bd:[ Li0>w0(16/48) Li1>w1(32/48) Ro0<w4(16/48) Ro1<w5(32/48) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output w4;    //: /sn:0 {0}(359,273)(359,337){1}
input w0;    //: /sn:0 {0}(356,147)(356,174){1}
//: {2}(358,176)(368,176)(368,223)(362,223)(362,252){3}
//: {4}(354,176)(261,176)(261,238){5}
input w1;    //: /sn:0 {0}(264,154)(264,164)(285,164)(285,212){1}
//: {2}(287,214)(357,214)(357,252){3}
//: {4}(283,214)(256,214)(256,238){5}
output w5;    //: /sn:0 {0}(258,259)(258,336){1}
//: enddecls

  //: joint g4 (w1) @(285, 214) /w:[ 2 1 4 -1 ]
  //: OUT g3 (w5) @(258,333) /sn:0 /R:3 /w:[ 1 ]
  //: OUT g2 (w4) @(359,334) /sn:0 /R:3 /w:[ 1 ]
  //: IN g1 (w1) @(264,152) /sn:0 /R:3 /w:[ 0 ]
  _GGXOR2 #(8) g6 (.I0(w0), .I1(w1), .Z(w4));   //: @(359,263) /sn:0 /R:3 /w:[ 3 3 0 ]
  //: joint g7 (w0) @(356, 176) /w:[ 2 1 4 -1 ]
  _GGAND2 #(6) g5 (.I0(w0), .I1(w1), .Z(w5));   //: @(258,249) /sn:0 /R:3 /w:[ 5 5 0 ]
  //: IN g0 (w0) @(356,145) /sn:0 /R:3 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin four_bit_adder
module four_bit_adder(w5, w3, w2, w1, w4, w0);
//: interface  /sz:(123, 80) /bd:[ Li0>w3(64/80) Li1>w2(48/80) Li2>w1(32/80) Li3>w0(16/80) Ro0<w5(32/80) Ro1<w4(16/80) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output w4;    //: /sn:0 {0}(304,462)(304,558)(324,558)(324,573){1}
input w3;    //: /sn:0 {0}(251,144)(251,346)(288,346)(288,361){1}
input w0;    //: /sn:0 {0}(449,146)(449,186)(402,186)(402,201){1}
input w1;    //: /sn:0 {0}(390,145)(390,186)(386,186)(386,201){1}
input w2;    //: /sn:0 {0}(320,147)(320,186)(370,186)(370,201){1}
output w5;    //: /sn:0 {0}(208,573)(208,600)(209,600)(209,615){1}
wire w7;    //: /sn:0 {0}(206,552)(206,333)(386,333)(386,314){1}
wire w12;    //: /sn:0 {0}(288,462)(288,537)(211,537)(211,552){1}
wire w8;    //: /sn:0 {0}(402,314)(402,350)(304,350)(304,361){1}
//: enddecls

  //: OUT g8 (w5) @(209,612) /sn:0 /R:3 /w:[ 1 ]
  full_adder g4 (.w8(w0), .w9(w1), .w10(w2), .w0(w8), .w1(w7));   //: @(354, 202) /sz:(64, 111) /R:3 /sn:0 /p:[ Ti0>1 Ti1>1 Ti2>1 Bo0<0 Bo1<1 ]
  //: IN g3 (w3) @(251,142) /sn:0 /R:3 /w:[ 0 ]
  //: IN g2 (w2) @(320,145) /sn:0 /R:3 /w:[ 0 ]
  //: IN g1 (w1) @(390,143) /sn:0 /R:3 /w:[ 0 ]
  _GGOR2 #(6) g6 (.I0(w12), .I1(w7), .Z(w5));   //: @(208,563) /sn:0 /R:3 /w:[ 1 0 0 ]
  //: OUT g7 (w4) @(324,570) /sn:0 /R:3 /w:[ 1 ]
  half_adder g5 (.w1(w3), .w0(w8), .w5(w12), .w4(w4));   //: @(272, 362) /sz:(48, 99) /R:3 /sn:0 /p:[ Ti0>1 Ti1>1 Bo0<0 Bo1<0 ]
  //: IN g0 (w0) @(449,144) /sn:0 /R:3 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin cross_two
module cross_two(w5, w3, w2, w1, w4, w0);
//: interface  /sz:(93, 80) /bd:[ Li0>w3(64/80) Li1>w2(48/80) Li2>w1(32/80) Li3>w0(16/80) Ro0<w5(32/80) Ro1<w4(16/80) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output w4;    //: /sn:0 {0}(440,590)(440,570)(433,570)(433,529){1}
input w3;    //: /sn:0 {0}(259,166)(259,262)(453,262)(453,277){1}
input w0;    //: /sn:0 {0}(580,168)(580,259)(458,259)(458,277){1}
input w1;    //: /sn:0 {0}(522,170)(522,339)(373,339)(373,354){1}
input w2;    //: /sn:0 {0}(322,165)(322,339)(368,339)(368,354){1}
output w5;    //: /sn:0 {0}(417,529)(417,569)(370,569)(370,620){1}
wire w6;    //: /sn:0 {0}(455,298)(455,413)(433,413)(433,428){1}
wire w9;    //: /sn:0 {0}(370,375)(370,413)(417,413)(417,428){1}
//: enddecls

  //: OUT g8 (w5) @(370,617) /sn:0 /R:3 /w:[ 1 ]
  _GGAND2 #(6) g4 (.I0(w0), .I1(w3), .Z(w6));   //: @(455,288) /sn:0 /R:3 /w:[ 1 1 0 ]
  //: IN g3 (w3) @(259,164) /sn:0 /R:3 /w:[ 0 ]
  //: IN g2 (w2) @(322,163) /sn:0 /R:3 /w:[ 0 ]
  //: IN g1 (w1) @(522,168) /sn:0 /R:3 /w:[ 0 ]
  half_adder g6 (.w0(w6), .w1(w9), .w4(w4), .w5(w5));   //: @(401, 429) /sz:(48, 99) /R:3 /sn:0 /p:[ Ti0>1 Ti1>1 Bo0<1 Bo1<0 ]
  //: OUT g7 (w4) @(440,587) /sn:0 /R:3 /w:[ 0 ]
  _GGAND2 #(6) g5 (.I0(w1), .I1(w2), .Z(w9));   //: @(370,365) /sn:0 /R:3 /w:[ 1 1 0 ]
  //: IN g0 (w0) @(580,166) /sn:0 /R:3 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin cross_three
module cross_three(w4, w3, w2, w1, w6, w7, w5, w0);
//: interface  /sz:(105, 112) /bd:[ Li0>w5(96/112) Li1>w4(80/112) Li2>w3(64/112) Li3>w2(48/112) Li4>w1(32/112) Li5>w0(16/112) Ro0<w7(32/112) Ro1<w6(16/112) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output w6;    //: /sn:0 {0}(379,560)(379,541)(363,541)(363,507)(346,507)(346,459){1}
output w7;    //: /sn:0 {0}(318,515)(318,474)(330,474)(330,459){1}
input w4;    //: /sn:0 {0}(258,119)(258,229)(245,229)(245,244){1}
input w3;    //: /sn:0 {0}(309,154)(309,231)(351,231)(351,246){1}
input w0;    //: /sn:0 {0}(489,112)(489,228)(485,228)(485,243){1}
input w1;    //: /sn:0 {0}(443,159)(443,228)(480,228)(480,243){1}
input w2;    //: /sn:0 {0}(372,120)(372,231)(356,231)(356,246){1}
input w5;    //: /sn:0 {0}(230,163)(230,229)(240,229)(240,244){1}
wire w8;    //: /sn:0 {0}(482,264)(482,325)(346,325)(346,346){1}
wire w14;    //: /sn:0 {0}(242,265)(242,331)(314,331)(314,346){1}
wire w11;    //: /sn:0 {0}(330,346)(330,308)(353,308)(353,267){1}
//: enddecls

  _GGAND2 #(6) g8 (.I0(w4), .I1(w5), .Z(w14));   //: @(242,255) /sn:0 /R:3 /w:[ 1 1 0 ]
  //: IN g4 (w4) @(258,117) /sn:0 /R:3 /w:[ 0 ]
  //: IN g3 (w3) @(309,152) /sn:0 /R:3 /w:[ 0 ]
  //: IN g2 (w2) @(372,118) /sn:0 /R:3 /w:[ 0 ]
  //: IN g1 (w1) @(443,157) /sn:0 /R:3 /w:[ 0 ]
  //: OUT g10 (w6) @(379,557) /sn:0 /R:3 /w:[ 0 ]
  _GGAND2 #(6) g6 (.I0(w0), .I1(w1), .Z(w8));   //: @(482,254) /sn:0 /R:3 /w:[ 1 1 0 ]
  full_adder g9 (.w8(w8), .w9(w11), .w10(w14), .w0(w6), .w1(w7));   //: @(298, 347) /sz:(64, 111) /R:3 /sn:0 /p:[ Ti0>1 Ti1>0 Ti2>1 Bo0<1 Bo1<1 ]
  _GGAND2 #(6) g7 (.I0(w2), .I1(w3), .Z(w11));   //: @(353,257) /sn:0 /R:3 /w:[ 1 1 1 ]
  //: OUT g11 (w7) @(318,512) /sn:0 /R:3 /w:[ 0 ]
  //: IN g5 (w5) @(230,161) /sn:0 /R:3 /w:[ 0 ]
  //: IN g0 (w0) @(489,110) /sn:0 /R:3 /w:[ 0 ]

endmodule
//: /netlistEnd

//: /netlistBegin full_adder
module full_adder(w10, w9, w8, w1, w0);
//: interface  /sz:(111, 64) /bd:[ Li0>w10(48/64) Li1>w9(32/64) Li2>w8(16/64) Ro0<w1(32/64) Ro1<w0(16/64) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
output w0;    //: /sn:0 {0}(395,548)(395,489)(379,489)(379,427){1}
input w10;    //: /sn:0 {0}(431,129)(431,172){1}
output w1;    //: /sn:0 {0}(299,554)(299,516)(305,516)(305,501){1}
input w8;    //: /sn:0 {0}(362,130)(362,157)(415,157)(415,172){1}
input w9;    //: /sn:0 {0}(363,326)(363,312)(294,312)(294,134){1}
wire w3;    //: /sn:0 {0}(431,273)(431,310)(379,310)(379,326){1}
wire w11;    //: /sn:0 {0}(308,480)(308,469)(363,469)(363,427){1}
wire w5;    //: /sn:0 {0}(303,480)(303,290)(415,290)(415,273){1}
//: enddecls

  _GGOR2 #(6) g8 (.I0(w11), .I1(w5), .Z(w1));   //: @(305,491) /sn:0 /R:3 /w:[ 0 0 1 ]
  //: IN g4 (w10) @(431,127) /sn:0 /R:3 /w:[ 0 ]
  //: IN g3 (w9) @(294,132) /sn:0 /R:3 /w:[ 1 ]
  //: IN g2 (w8) @(362,128) /sn:0 /R:3 /w:[ 0 ]
  half_adder g1 (.w1(w9), .w0(w3), .w5(w11), .w4(w0));   //: @(347, 327) /sz:(48, 99) /R:3 /sn:0 /p:[ Ti0>0 Ti1>1 Bo0<1 Bo1<1 ]
  //: OUT g6 (w1) @(299,551) /sn:0 /R:3 /w:[ 0 ]
  //: OUT g5 (w0) @(395,545) /sn:0 /R:3 /w:[ 0 ]
  half_adder g0 (.w1(w8), .w0(w10), .w5(w5), .w4(w3));   //: @(399, 173) /sz:(48, 99) /R:3 /sn:0 /p:[ Ti0>1 Ti1>1 Bo0<1 Bo1<0 ]

endmodule
//: /netlistEnd

//: /netlistBegin cross_four
module cross_four(w4, w3, w2, w1, w6, w7, w9, w5, w0, w8);
//: interface  /sz:(99, 144) /bd:[ Li0>w7(128/144) Li1>w6(112/144) Li2>w5(96/144) Li3>w4(80/144) Li4>w3(64/144) Li5>w2(48/144) Li6>w1(32/144) Li7>w0(16/144) Ro0<w9(32/144) Ro1<w8(16/144) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input w6;    //: /sn:0 {0}(113,108)(113,162)(138,162)(138,177){1}
input w7;    //: /sn:0 {0}(154,108)(154,162)(143,162)(143,177){1}
input w4;    //: /sn:0 {0}(214,94)(214,156)(230,156)(230,171){1}
input w3;    //: /sn:0 {0}(357,93)(357,154)(341,154)(341,169){1}
input w0;    //: /sn:0 {0}(462,108)(462,169)(443,169)(443,184){1}
input w1;    //: /sn:0 {0}(421,108)(421,169)(438,169)(438,184){1}
output w8;    //: /sn:0 {0}(308,401)(308,462)(337,462)(337,477){1}
input w2;    //: /sn:0 {0}(316,93)(316,154)(336,154)(336,169){1}
input w5;    //: /sn:0 {0}(255,94)(255,156)(235,156)(235,171){1}
output w9;    //: /sn:0 {0}(292,401)(292,465)(275,465)(275,480){1}
wire w16;    //: /sn:0 {0}(276,276)(276,235)(232,235)(232,192){1}
wire w13;    //: /sn:0 {0}(292,276)(292,205)(338,205)(338,190){1}
wire w19;    //: /sn:0 {0}(140,198)(140,249)(260,249)(260,276){1}
wire w10;    //: /sn:0 {0}(308,276)(308,260)(440,260)(440,205){1}
//: enddecls

  _GGAND2 #(6) g8 (.I0(w0), .I1(w1), .Z(w10));   //: @(440,195) /sn:0 /R:3 /w:[ 1 1 1 ]
  //: IN g4 (w4) @(214,92) /sn:0 /R:3 /w:[ 0 ]
  //: IN g3 (w3) @(357,91) /sn:0 /R:3 /w:[ 0 ]
  //: IN g2 (w2) @(316,91) /sn:0 /R:3 /w:[ 0 ]
  //: IN g1 (w1) @(421,106) /sn:0 /R:3 /w:[ 0 ]
  _GGAND2 #(6) g10 (.I0(w5), .I1(w4), .Z(w16));   //: @(232,182) /sn:0 /R:3 /w:[ 1 1 1 ]
  //: IN g6 (w6) @(113,106) /sn:0 /R:3 /w:[ 0 ]
  _GGAND2 #(6) g9 (.I0(w3), .I1(w2), .Z(w13));   //: @(338,180) /sn:0 /R:3 /w:[ 1 1 1 ]
  //: IN g7 (w7) @(154,106) /sn:0 /R:3 /w:[ 0 ]
  four_bit_adder g12 (.w0(w10), .w1(w13), .w2(w16), .w3(w19), .w4(w8), .w5(w9));   //: @(244, 277) /sz:(80, 123) /R:3 /sn:0 /p:[ Ti0>0 Ti1>0 Ti2>0 Ti3>1 Bo0<0 Bo1<0 ]
  //: OUT g14 (w9) @(275,477) /sn:0 /R:3 /w:[ 1 ]
  _GGAND2 #(6) g11 (.I0(w7), .I1(w6), .Z(w19));   //: @(140,188) /sn:0 /R:3 /w:[ 1 1 0 ]
  //: IN g5 (w5) @(255,92) /sn:0 /R:3 /w:[ 0 ]
  //: IN g0 (w0) @(462,106) /sn:0 /R:3 /w:[ 0 ]
  //: OUT g13 (w8) @(337,474) /sn:0 /R:3 /w:[ 1 ]

endmodule
//: /netlistEnd

