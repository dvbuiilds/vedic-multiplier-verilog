//: version "2.1"
//: property encoding = "utf-8"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "FLIPFLOP.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg w0;    //: /sn:0 {0}(126,124)(149,124){1}
//: {2}(153,124)(202,124)(202,158)(230,158){3}
//: {4}(151,126)(151,300)(170,300){5}
wire w6;    //: /sn:0 {0}(358,180)(375,180){1}
//: {2}(379,180)(433,180){3}
//: {4}(377,182)(377,264)(320,264)(320,279)(330,279){5}
wire w7;    //: /sn:0 {0}(330,284)(316,284)(316,290)(248,290){1}
wire w4;    //: /sn:0 {0}(337,177)(328,177)(328,144)(261,144)(261,161)(251,161){1}
wire w3;    //: /sn:0 {0}(115,224)(215,224){1}
//: {2}(217,222)(217,163)(230,163){3}
//: {4}(217,226)(217,287)(227,287){5}
wire w8;    //: /sn:0 {0}(186,300)(217,300)(217,292)(227,292){1}
wire w5;    //: /sn:0 {0}(351,282)(382,282){1}
//: {2}(386,282)(422,282)(422,281)(437,281){3}
//: {4}(384,280)(384,197)(327,197)(327,182)(337,182){5}
//: enddecls

  _GGNOR2 #(4) g4 (.I0(w4), .I1(w5), .Z(w6));   //: @(348,180) /sn:0 /w:[ 0 5 0 ]
  _GGCLOCK_P20_0_50 g8 (.Z(w3));   //: @(102,224) /sn:0 /w:[ 0 ] /omega:20 /phi:0 /duty:50
  //: comment g16 @(319,311) /sn:0
  //: /line:"R"
  //: /end
  _GGNAND2 #(4) g3 (.I0(w0), .I1(w3), .Z(w4));   //: @(241,161) /sn:0 /w:[ 3 3 1 ]
  _GGNAND2 #(4) g2 (.I0(w3), .I1(w8), .Z(w7));   //: @(238,290) /sn:0 /w:[ 5 1 1 ]
  //: joint g1 (w3) @(217, 224) /w:[ -1 2 1 4 ]
  //: LED g10 (w6) @(440,180) /sn:0 /R:3 /w:[ 3 ] /type:0
  //: joint g6 (w6) @(377, 180) /w:[ 2 -1 1 4 ]
  //: joint g9 (w0) @(151, 124) /w:[ 2 -1 1 4 ]
  //: joint g7 (w5) @(384, 282) /w:[ 2 4 1 -1 ]
  //: comment g12 @(63,118) /sn:0
  //: /line:"D"
  //: /end
  _GGNOR2 #(4) g5 (.I0(w6), .I1(w7), .Z(w5));   //: @(341,282) /sn:0 /w:[ 5 0 0 ]
  //: LED g11 (w5) @(444,281) /sn:0 /R:3 /w:[ 3 ] /type:0
  //: comment g14 @(53,221) /sn:0
  //: /line:"CP"
  //: /end
  _GGNBUF #(2) g15 (.I(w0), .Z(w8));   //: @(176,300) /sn:0 /w:[ 5 0 ]
  //: SWITCH g0 (w0) @(109,124) /sn:0 /w:[ 0 ] /st:1 /dn:1
  //: comment g13 @(308,122) /sn:0
  //: /line:"S"
  //: /end

endmodule
//: /netlistEnd

