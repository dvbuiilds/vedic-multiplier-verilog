//: version "2.1"
//: property encoding = "utf-8"
//: property locale = "en"
//: property prefix = "_GG"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg w3;    //: /sn:0 {0}(92,348)(178,348)(178,347)(193,347){1}
reg w0;    //: /sn:0 {0}(90,100)(154,100){1}
//: {2}(158,100)(260,100){3}
//: {4}(156,102)(156,176)(189,176){5}
reg w1;    //: /sn:0 {0}(92,183)(155,183){1}
//: {2}(159,183)(176,183)(176,181)(189,181){3}
//: {4}(157,185)(157,260)(190,260){5}
reg w2;    //: /sn:0 {0}(94,265)(155,265){1}
//: {2}(159,265)(190,265){3}
//: {4}(157,267)(157,342)(193,342){5}
wire w6;    //: /sn:0 {0}(261,179)(210,179){1}
wire w12;    //: /sn:0 {0}(214,345)(268,345){1}
wire w9;    //: /sn:0 {0}(211,263)(265,263){1}
//: enddecls

  //: joint g8 (w1) @(157, 183) /w:[ 2 -1 1 4 ]
  _GGXOR2 #(8) g4 (.I0(w0), .I1(w1), .Z(w6));   //: @(200,179) /sn:0 /w:[ 5 3 1 ]
  //: SWITCH g3 (w3) @(75,348) /sn:0 /w:[ 0 ] /st:1 /dn:1
  //: SWITCH g2 (w2) @(77,265) /sn:0 /w:[ 0 ] /st:1 /dn:1
  //: SWITCH g1 (w1) @(75,183) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: LED g10 (w0) @(267,100) /sn:0 /R:3 /w:[ 3 ] /type:0
  _GGXOR2 #(8) g6 (.I0(w2), .I1(w3), .Z(w12));   //: @(204,345) /sn:0 /w:[ 5 1 0 ]
  //: joint g9 (w2) @(157, 265) /w:[ 2 -1 1 4 ]
  //: joint g7 (w0) @(156, 100) /w:[ 2 -1 1 4 ]
  //: LED g12 (w9) @(272,263) /sn:0 /R:3 /w:[ 1 ] /type:0
  //: LED g11 (w6) @(268,179) /sn:0 /R:3 /w:[ 0 ] /type:0
  _GGXOR2 #(8) g5 (.I0(w1), .I1(w2), .Z(w9));   //: @(201,263) /sn:0 /w:[ 5 3 0 ]
  //: SWITCH g0 (w0) @(73,100) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: LED g13 (w12) @(275,345) /sn:0 /R:3 /w:[ 1 ] /type:0

endmodule
//: /netlistEnd

