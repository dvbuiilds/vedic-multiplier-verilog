//: version "2.1"
//: property encoding = "utf-8"
//: property locale = "en"
//: property prefix = "_GG"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg w3;    //: /sn:0 {0}(106,100)(282,100)(282,102)(292,102){1}
//: {2}(294,100)(294,91)(367,91)(367,158)(380,158){3}
//: {4}(294,104)(294,222)(318,222){5}
reg w1;    //: /sn:0 {0}(105,167)(166,167){1}
//: {2}(170,167)(189,167)(189,189)(202,189){3}
//: {4}(168,169)(168,258)(215,258){5}
reg w2;    //: /sn:0 {0}(107,248)(126,248){1}
//: {2}(130,248)(189,248)(189,194)(202,194){3}
//: {4}(128,250)(128,270)(146,270){5}
wire w7;    //: /sn:0 {0}(284,228)(303,228)(303,227)(318,227){1}
wire w4;    //: /sn:0 {0}(162,270)(200,270)(200,263)(215,263){1}
wire w8;    //: /sn:0 {0}(401,161)(420,161)(420,160)(435,160){1}
wire w17;    //: /sn:0 {0}(401,238)(435,238){1}
wire w14;    //: /sn:0 {0}(339,225)(365,225)(365,235)(380,235){1}
wire w11;    //: /sn:0 {0}(236,261)(365,261)(365,240)(380,240){1}
wire w5;    //: /sn:0 {0}(223,192)(248,192){1}
//: {2}(252,192)(367,192)(367,163)(380,163){3}
//: {4}(250,194)(250,228)(268,228){5}
//: enddecls

  _GGAND2 #(6) g8 (.I0(w3), .I1(w7), .Z(w14));   //: @(329,225) /sn:0 /w:[ 5 1 0 ]
  _GGXOR2 #(8) g4 (.I0(w3), .I1(w5), .Z(w8));   //: @(391,161) /sn:0 /w:[ 3 3 0 ]
  _GGXOR2 #(8) g3 (.I0(w1), .I1(w2), .Z(w5));   //: @(213,192) /sn:0 /w:[ 3 3 0 ]
  //: SWITCH g2 (w2) @(90,248) /sn:0 /w:[ 0 ] /st:1 /dn:1
  //: SWITCH g1 (w1) @(88,167) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: joint g10 (w2) @(128, 248) /w:[ 2 -1 1 4 ]
  _GGNBUF #(2) g6 (.I(w5), .Z(w7));   //: @(274,228) /sn:0 /w:[ 5 0 ]
  _GGOR2 #(6) g9 (.I0(w14), .I1(w11), .Z(w17));   //: @(391,238) /sn:0 /w:[ 1 1 0 ]
  _GGAND2 #(6) g7 (.I0(w1), .I1(w4), .Z(w11));   //: @(226,261) /sn:0 /w:[ 5 1 0 ]
  //: joint g12 (w5) @(250, 192) /w:[ 2 -1 1 4 ]
  //: LED g14 (w8) @(442,160) /sn:0 /R:3 /w:[ 1 ] /type:0
  //: joint g11 (w1) @(168, 167) /w:[ 2 -1 1 4 ]
  _GGNBUF #(2) g5 (.I(w2), .Z(w4));   //: @(152,270) /sn:0 /w:[ 5 0 ]
  //: SWITCH g0 (w3) @(89,100) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: LED g15 (w17) @(442,238) /sn:0 /R:3 /w:[ 1 ] /type:0
  //: joint g13 (w3) @(294, 102) /w:[ -1 2 1 4 ]

endmodule
//: /netlistEnd

