//: version "2.1"
//: property encoding = "utf-8"
//: property locale = "en"
//: property prefix = "_GG"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg w2;    //: /sn:0 {0}(45,153)(59,153)(59,150){1}
//: {2}(61,148)(73,148)(73,150)(158,150){3}
//: {4}(59,146)(59,99)(80,99){5}
wire w13;    //: /sn:0 {0}(271,95)(252,95)(252,96){1}
//: {2}(254,98)(263,98)(263,100)(271,100){3}
//: {4}(250,98)(245,98){5}
wire w7;    //: /sn:0 {0}(177,67)(209,67)(209,95)(224,95){1}
wire w4;    //: /sn:0 {0}(101,97)(139,97){1}
//: {2}(141,95)(141,69)(156,69){3}
//: {4}(141,99)(141,145)(158,145){5}
wire w0;    //: /sn:0 {0}(80,94)(55,94)(55,66){1}
//: {2}(57,64)(156,64){3}
//: {4}(55,62)(55,34)(40,34){5}
wire w10;    //: /sn:0 {0}(224,100)(194,100)(194,148)(179,148){1}
wire w1;    //: /sn:0 {0}(317,97)(307,97)(307,98)(292,98){1}
//: enddecls

  //: joint g8 (w0) @(55, 64) /w:[ 2 4 -1 1 ]
  _GGNAND2 #(4) g4 (.I0(w4), .I1(w2), .Z(w10));   //: @(169,148) /sn:0 /w:[ 5 3 1 ]
  _GGNAND2 #(4) g3 (.I0(w0), .I1(w4), .Z(w7));   //: @(167,67) /sn:0 /w:[ 3 3 0 ]
  _GGNAND2 #(4) g2 (.I0(w0), .I1(w2), .Z(w4));   //: @(91,97) /sn:0 /w:[ 0 5 0 ]
  //: SWITCH g1 (w2) @(28,153) /sn:0 /w:[ 0 ] /st:0 /dn:1
  _GGNAND2 #(4) g10 (.I0(w13), .I1(w13), .Z(w1));   //: @(282,98) /sn:0 /w:[ 0 3 1 ]
  //: LED g6 (w1) @(324,97) /sn:0 /R:3 /w:[ 0 ] /type:0
  //: joint g9 (w2) @(59, 148) /w:[ 2 4 -1 1 ]
  //: joint g7 (w4) @(141, 97) /w:[ -1 2 1 4 ]
  //: joint g11 (w13) @(252, 98) /w:[ 2 1 4 -1 ]
  _GGNAND2 #(4) g5 (.I0(w7), .I1(w10), .Z(w13));   //: @(235,98) /sn:0 /w:[ 1 0 5 ]
  _GGCLOCK_P100_0_50 g0 (.Z(w0));   //: @(27,34) /sn:0 /w:[ 5 ] /omega:100 /phi:0 /duty:50

endmodule
//: /netlistEnd

