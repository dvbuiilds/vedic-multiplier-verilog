//: version "2.1"
//: property encoding = "utf-8"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "GREYCODE.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg w0;    //: /sn:0 {0}(332,425)(332,458)(254,458){1}
//: {2}(252,456)(252,383)(254,383)(254,329){3}
//: {4}(252,460)(252,541){5}
reg w3;    //: /sn:0 {0}(498,437)(498,471)(500,471)(500,539){1}
reg w1;    //: /sn:0 {0}(339,539)(339,459){1}
//: {2}(341,457)(407,457)(407,429){3}
//: {4}(339,455)(339,441)(337,441)(337,425){5}
reg w2;    //: /sn:0 {0}(412,429)(412,456){1}
//: {2}(414,458)(493,458)(493,437){3}
//: {4}(412,460)(412,479)(417,479)(417,537){5}
wire w13;    //: /sn:0 {0}(410,326)(410,408){1}
wire w4;    //: /sn:0 {0}(335,328)(335,404){1}
wire w5;    //: /sn:0 {0}(496,416)(496,387)(497,387)(497,327){1}
//: enddecls

  //: joint g4 (w0) @(252, 458) /w:[ 1 2 -1 4 ]
  _GGXOR2 #(8) g16 (.I0(w1), .I1(w2), .Z(w13));   //: @(410,418) /sn:0 /R:1 /w:[ 3 0 1 ]
  //: SWITCH g3 (w3) @(500,553) /sn:0 /R:1 /w:[ 1 ] /st:0 /dn:1
  //: LED g17 (w4) @(335,321) /sn:0 /w:[ 0 ] /type:0
  //: SWITCH g2 (w2) @(417,551) /sn:0 /R:1 /w:[ 5 ] /st:0 /dn:1
  //: SWITCH g1 (w1) @(339,553) /sn:0 /R:1 /w:[ 0 ] /st:0 /dn:1
  //: LED g18 (w0) @(254,322) /sn:0 /w:[ 3 ] /type:0
  _GGXOR2 #(8) g10 (.I0(w0), .I1(w1), .Z(w4));   //: @(335,414) /sn:0 /R:1 /w:[ 0 5 1 ]
  //: joint g6 (w2) @(412, 458) /w:[ 2 1 -1 4 ]
  //: joint g5 (w1) @(339, 457) /w:[ 2 4 -1 1 ]
  _GGXOR2 #(8) g14 (.I0(w2), .I1(w3), .Z(w5));   //: @(496,426) /sn:0 /R:1 /w:[ 3 0 0 ]
  //: LED g15 (w13) @(410,319) /sn:0 /w:[ 0 ] /type:0
  //: SWITCH g0 (w0) @(252,555) /sn:0 /R:1 /w:[ 5 ] /st:0 /dn:1
  //: LED g13 (w5) @(497,320) /sn:0 /w:[ 1 ] /type:0

endmodule
//: /netlistEnd

