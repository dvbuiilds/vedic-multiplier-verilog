//: version "2.1"
//: property encoding = "utf-8"
//: property locale = "en"
//: property prefix = "_GG"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg w0;    //: /sn:0 {0}(90,45)(106,45){1}
//: {2}(110,45)(117,45)(117,66)(130,66){3}
//: {4}(108,47)(108,212)(183,212){5}
reg w1;    //: /sn:0 {0}(91,92)(95,92){1}
//: {2}(99,92)(117,92)(117,71)(130,71){3}
//: {4}(97,94)(97,217)(183,217){5}
wire w13;    //: /sn:0 {0}(316,191)(308,191)(308,193)(258,193){1}
wire w6;    //: /sn:0 {0}(235,104)(205,104){1}
wire w7;    //: /sn:0 {0}(237,190)(218,190)(218,170)(203,170){1}
wire w10;    //: /sn:0 {0}(237,195)(219,195)(219,215)(204,215){1}
wire w2;    //: /sn:0 {0}(86,129)(168,129){1}
//: {2}(170,127)(170,106)(184,106){3}
//: {4}(170,131)(170,167)(182,167){5}
wire w5;    //: /sn:0 {0}(151,69)(155,69){1}
//: {2}(159,69)(171,69)(171,101)(184,101){3}
//: {4}(157,71)(157,172)(182,172){5}
//: enddecls

  //: joint g8 (w2) @(170, 129) /w:[ -1 2 1 4 ]
  _GGXOR2 #(8) g4 (.I0(w5), .I1(w2), .Z(w6));   //: @(195,104) /sn:0 /w:[ 3 3 1 ]
  //: comment g16 @(27,88) /sn:0
  //: /line:"  B"
  //: /end
  _GGXOR2 #(8) g3 (.I0(w0), .I1(w1), .Z(w5));   //: @(141,69) /sn:0 /w:[ 3 3 0 ]
  //: comment g17 @(261,102) /sn:0
  //: /line:"SUM"
  //: /end
  _GGCLOCK_P50_0_50 g2 (.Z(w2));   //: @(73,129) /sn:0 /w:[ 0 ] /omega:50 /phi:0 /duty:50
  //: SWITCH g1 (w1) @(74,92) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: comment g18 @(334,186) /sn:0
  //: /line:"C OUT"
  //: /end
  //: joint g10 (w0) @(108, 45) /w:[ 2 -1 1 4 ]
  _GGAND2 #(6) g6 (.I0(w0), .I1(w1), .Z(w10));   //: @(194,215) /sn:0 /w:[ 5 5 1 ]
  //: joint g9 (w5) @(157, 69) /w:[ 2 -1 1 4 ]
  _GGOR2 #(6) g7 (.I0(w7), .I1(w10), .Z(w13));   //: @(248,193) /sn:0 /w:[ 0 0 1 ]
  //: LED g12 (w6) @(242,104) /sn:0 /R:3 /w:[ 0 ] /type:0
  //: comment g14 @(22,123) /sn:0
  //: /line:"C IN"
  //: /end
  //: joint g11 (w1) @(97, 92) /w:[ 2 -1 1 4 ]
  _GGAND2 #(6) g5 (.I0(w2), .I1(w5), .Z(w7));   //: @(193,170) /sn:0 /w:[ 5 5 1 ]
  //: comment g15 @(27,35) /sn:0
  //: /line:"  A"
  //: /end
  //: SWITCH g0 (w0) @(73,45) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: LED g13 (w13) @(323,191) /sn:0 /R:3 /w:[ 0 ] /type:0

endmodule
//: /netlistEnd

