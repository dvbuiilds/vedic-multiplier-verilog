//: version "2.1"
//: property encoding = "utf-8"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "1:4-DEMUX.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg w0;    //: /sn:0 {0}(181,221)(499,221){1}
//: {2}(503,221)(513,221)(513,222)(548,222){3}
//: {4}(501,223)(501,328){5}
//: {6}(503,330)(547,330){7}
//: {8}(501,332)(501,441){9}
//: {10}(503,443)(550,443){11}
//: {12}(501,445)(501,553)(551,553){13}
reg w30;    //: /sn:0 {0}(350,80)(350,96){1}
//: {2}(352,98)(424,98)(424,109){3}
//: {4}(350,100)(350,273){5}
//: {6}(352,275)(362,275)(362,276)(547,276){7}
//: {8}(350,277)(350,499)(551,499){9}
reg w29;    //: /sn:0 {0}(265,79)(265,110){1}
//: {2}(267,112)(366,112)(366,129){3}
//: {4}(265,114)(265,402){5}
//: {6}(267,404)(277,404)(277,407)(550,407){7}
//: {8}(265,406)(265,517)(551,517){9}
reg w1;    //: /sn:0 {0}(548,204)(483,204)(483,311){1}
//: {2}(485,313)(495,313)(495,312)(547,312){3}
//: {4}(483,315)(483,422){5}
//: {6}(485,424)(495,424)(495,425)(550,425){7}
//: {8}(483,426)(483,531){9}
//: {10}(485,533)(495,533)(495,535)(551,535){11}
//: {12}(483,535)(483,544)(176,544){13}
wire w6;    //: /sn:0 {0}(424,125)(424,166){1}
//: {2}(426,168)(548,168){3}
//: {4}(424,170)(424,389)(550,389){5}
wire w7;    //: /sn:0 {0}(773,167)(778,167){1}
//: {2}(782,167)(796,167)(796,166)(800,166){3}
//: {4}(780,165)(780,168)(744,168){5}
wire w22;    //: /sn:0 {0}(747,499)(780,499)(780,500)(795,500){1}
wire w12;    //: /sn:0 {0}(743,276)(796,276)(796,293)(811,293){1}
wire w17;    //: /sn:0 {0}(746,389)(784,389)(784,413)(799,413){1}
wire w5;    //: /sn:0 {0}(366,145)(366,184){1}
//: {2}(368,186)(548,186){3}
//: {4}(366,188)(366,294)(547,294){5}
//: enddecls

  //: SWITCH g8 (w1) @(159,544) /sn:0 /w:[ 13 ] /st:0 /dn:1
  four_input_and_gate g4 (.iNPUT1(w30), .INPUT2(w29), .INPUT3(w1), .INPUT4(w0), .OUTPUT1(w22));   //: @(552, 481) /sz:(194, 90) /sn:0 /p:[ Li0>9 Li1>9 Li2>11 Li3>13 Ro0<0 ]
  //: joint g16 (w1) @(483, 533) /w:[ 10 9 -1 12 ]
  four_input_and_gate g3 (.iNPUT1(w6), .INPUT2(w29), .INPUT3(w1), .INPUT4(w0), .OUTPUT1(w17));   //: @(551, 371) /sz:(194, 90) /sn:0 /p:[ Li0>5 Li1>7 Li2>7 Li3>11 Ro0<0 ]
  //: LED g26 (w17) @(806,413) /sn:0 /R:3 /w:[ 1 ] /type:0
  //: joint g17 (w30) @(350, 98) /w:[ 2 1 -1 4 ]
  four_input_and_gate g2 (.iNPUT1(w30), .INPUT2(w5), .INPUT3(w1), .INPUT4(w0), .OUTPUT1(w12));   //: @(548, 258) /sz:(194, 90) /sn:0 /p:[ Li0>7 Li1>5 Li2>3 Li3>7 Ro0<0 ]
  //: joint g23 (w29) @(265, 404) /w:[ 6 5 -1 8 ]
  //: LED g24 (w7) @(807,166) /sn:0 /R:3 /w:[ 3 ] /type:0
  four_input_and_gate g1 (.iNPUT1(w6), .INPUT2(w5), .INPUT3(w1), .INPUT4(w0), .OUTPUT1(w7));   //: @(549, 150) /sz:(194, 90) /sn:0 /p:[ Li0>3 Li1>3 Li2>0 Li3>3 Ro0<5 ]
  //: joint g18 (w30) @(350, 275) /w:[ 6 5 -1 8 ]
  //: LED g25 (w12) @(818,293) /sn:0 /R:3 /w:[ 1 ] /type:0
  _GGNBUF #(2) g10 (.I(w29), .Z(w5));   //: @(366,135) /sn:0 /R:3 /w:[ 3 0 ]
  //: joint g6 (w0) @(501, 330) /w:[ 6 5 -1 8 ]
  //: joint g7 (w0) @(501, 443) /w:[ 10 9 -1 12 ]
  _GGNBUF #(2) g9 (.I(w30), .Z(w6));   //: @(424,115) /sn:0 /R:3 /w:[ 3 0 ]
  //: joint g22 (w6) @(424, 168) /w:[ 2 1 -1 4 ]
  //: SWITCH g12 (w30) @(350,67) /sn:0 /R:3 /w:[ 0 ] /st:0 /dn:1
  //: joint g28 (w7) @(780, 167) /w:[ 2 -1 1 4 ]
  //: joint g14 (w1) @(483, 313) /w:[ 2 1 -1 4 ]
  //: joint g5 (w0) @(501, 221) /w:[ 2 -1 1 4 ]
  //: SWITCH g11 (w29) @(265,66) /sn:0 /R:3 /w:[ 0 ] /st:0 /dn:1
  //: joint g21 (w5) @(366, 186) /w:[ 2 1 -1 4 ]
  //: comment g19 @(249,17) /sn:0
  //: /line:"S1"
  //: /end
  //: comment g20 @(336,17) /sn:0
  //: /line:"S0"
  //: /end
  //: joint g15 (w1) @(483, 424) /w:[ 6 5 -1 8 ]
  //: SWITCH g0 (w0) @(164,221) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: LED g27 (w22) @(802,500) /sn:0 /R:3 /w:[ 1 ] /type:0
  //: joint g13 (w29) @(265, 112) /w:[ 2 1 -1 4 ]

endmodule
//: /netlistEnd

//: /netlistBegin four_input_and_gate
module four_input_and_gate(INPUT3, INPUT2, iNPUT1, INPUT4, OUTPUT1);
//: interface  /sz:(194, 90) /bd:[ Li0>INPUT4(64/80) Li1>INPUT3(48/80) Li2>INPUT2(32/80) Li3>iNPUT1(16/80) Ro0<OUTPUT1(16/80) ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
input iNPUT1;    //: {0}(93,45)(50:132,45)(132,65)(147,65){1}
output OUTPUT1;    //: /sn:0 {0}(436,100)(352,100)(352,134)(287,134){1}
input INPUT4;    //: /sn:0 {0}(95,136)(266,136){1}
input INPUT3;    //: /sn:0 {0}(95,104)(207,104){1}
input INPUT2;    //: {0}(95,73)(50:132,73)(132,70)(147,70){1}
wire w0;    //: /sn:0 {0}(228,102)(251,102)(251,131)(266,131){1}
wire w2;    //: /sn:0 {0}(168,68)(191,68)(191,99)(207,99){1}
//: enddecls

  //: IN g4 (INPUT3) @(93,104) /sn:0 /w:[ 0 ]
  //: IN g3 (INPUT2) @(93,73) /sn:0 /w:[ 0 ]
  //: IN g2 (iNPUT1) @(91,45) /sn:0 /w:[ 0 ]
  _GGAND2 #(6) g1 (.I0(w2), .I1(INPUT3), .Z(w0));   //: @(218,102) /sn:0 /w:[ 1 1 0 ]
  _GGAND2 #(6) g6 (.I0(w0), .I1(INPUT4), .Z(OUTPUT1));   //: @(277,134) /sn:0 /w:[ 1 1 1 ]
  //: IN g7 (INPUT4) @(93,136) /sn:0 /w:[ 0 ]
  //: OUT g5 (OUTPUT1) @(433,100) /sn:0 /w:[ 0 ]
  _GGAND2 #(6) g0 (.I0(iNPUT1), .I1(INPUT2), .Z(w2));   //: @(158,68) /sn:0 /w:[ 1 1 0 ]

endmodule
//: /netlistEnd

