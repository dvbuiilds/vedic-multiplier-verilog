//: version "2.1"
//: property encoding = "utf-8"
//: property locale = "en"
//: property prefix = "_GG"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg w1;    //: /sn:0 {0}(128,112)(74,112)(74,157){1}
//: {2}(72,159)(59,159){3}
//: {4}(74,161)(74,199)(238,199){5}
wire w13;    //: /sn:0 {0}(393,112)(425,112)(425,110)(436,110){1}
wire w7;    //: /sn:0 {0}(321,109)(282,109)(282,49)(255,49){1}
wire w4;    //: /sn:0 {0}(149,110)(217,110){1}
//: {2}(221,110)(227,110)(227,194)(238,194){3}
//: {4}(219,108)(219,51)(234,51){5}
wire w0;    //: /sn:0 {0}(128,107)(67,107)(67,62){1}
//: {2}(67,58)(67,46)(234,46){3}
//: {4}(65,60)(52,60){5}
wire w10;    //: /sn:0 {0}(321,114)(274,114)(274,197)(259,197){1}
wire w2;    //: /sn:0 {0}(372,109)(354,109){1}
//: {2}(350,109)(346,109)(346,112)(342,112){3}
//: {4}(352,111)(352,114)(372,114){5}
//: enddecls

  //: joint g8 (w1) @(74, 159) /w:[ -1 1 2 4 ]
  _GGNOR2 #(4) g4 (.I0(w4), .I1(w1), .Z(w10));   //: @(249,197) /sn:0 /w:[ 3 5 1 ]
  _GGNOR2 #(4) g3 (.I0(w0), .I1(w4), .Z(w7));   //: @(245,49) /sn:0 /w:[ 3 5 1 ]
  _GGNOR2 #(4) g2 (.I0(w0), .I1(w1), .Z(w4));   //: @(139,110) /sn:0 /w:[ 0 0 0 ]
  //: SWITCH g1 (w1) @(42,159) /sn:0 /w:[ 3 ] /st:0 /dn:1
  _GGNOR2 #(4) g10 (.I0(w2), .I1(w2), .Z(w13));   //: @(383,112) /sn:0 /w:[ 0 5 0 ]
  //: joint g6 (w4) @(219, 110) /w:[ 2 4 1 -1 ]
  //: LED g9 (w13) @(443,110) /sn:0 /R:3 /w:[ 1 ] /type:0
  //: joint g7 (w0) @(67, 60) /w:[ -1 2 4 1 ]
  //: joint g11 (w2) @(352, 109) /w:[ 1 -1 2 4 ]
  _GGNOR2 #(4) g5 (.I0(w7), .I1(w10), .Z(w2));   //: @(332,112) /sn:0 /w:[ 0 0 3 ]
  _GGCLOCK_P100_0_50 g0 (.Z(w0));   //: @(39,60) /sn:0 /w:[ 5 ] /omega:100 /phi:0 /duty:50

endmodule
//: /netlistEnd

